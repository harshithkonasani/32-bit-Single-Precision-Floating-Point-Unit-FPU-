`timescale 1ns / 1ps

module fpu_division(
    input [31:0] float_num1,
    input [31:0] float_num2,
    output reg [31:0] div_result,
    output [7:0]pos,
    output [7:0] exponent1, exponent2,
    output [22:0] mantissa1, mantissa2,
    output sign1, sign2
);

// Partition of floating-point numbers
wire [7:0] exp_num1, exp_num2;
wire [23:0] mantissa_num1, mantissa_num2;
wire sign_num1, sign_num2;

// Outputs from various components
wire [7:0] exponent_subtract;
wire [7:0] adjusted_exponent;
reg sign_out;

wire exception;

// Normalizer outputs
reg [7:0] normalized_exponent = 8'b0;  // Initialize to avoid unset bits
reg [23:0] normalized_mantissa = 24'b0;  // Initialize to avoid unset bits

// Assign input partitions 
assign sign_num1 = float_num1[31];
assign exp_num1 = float_num1[30:23];
assign sign_num2 = float_num2[31];
assign exp_num2 = float_num2[30:23];

// Check for division by zero
assign exception = (float_num2 == 32'b0) ? 1'b1 : 1'b0;

// Ensure mantissa is set correctly
assign mantissa_num1 = (exception) ? 24'b0 : {1'b1, float_num1[22:0]};
assign mantissa_num2 = (exception) ? 24'b0 : {1'b1, float_num2[22:0]};

assign exponent1 = exp_num1;
assign exponent2 = exp_num2;
assign sign1 = sign_num1;
assign sign2 = sign_num2;
assign mantissa1 = mantissa_num1;
assign mantissa2 = mantissa_num2;

// Exponent difference calculation
assign exponent_subtract = exp_num1 - exp_num2;  // Direct subtraction

// Adjust the exponent (bias correction of 127)
assign adjusted_exponent = exponent_subtract[7:0] + 8'b01111111;  // Keep only 8 bits

// Mantissa division result (48-bit precision)
reg [47:0] mantissa_div_result;  
reg [7:0] position;  // 6-bit position
reg [47:0] shifted_mantissa;  

//intermediate division result
wire [47:0] intermediate_div_result;  

divider d0(.mantissa_num1(mantissa_num1),.mantissa_num2(mantissa_num2),.mantissa_div_result(intermediate_div_result));

always @(*) begin
    if (exception) begin
        mantissa_div_result = 48'b0; // Set to zero if division by zero occurs
    end else begin
        mantissa_div_result = intermediate_div_result;
    end

    case (mantissa_div_result)
        48'b1??????????????????????????????????????????????? : position = 8'd0;
        48'b01?????????????????????????????????????????????? : position = 8'd1;
        48'b001????????????????????????????????????????????? : position = 8'd2;
        48'b0001???????????????????????????????????????????? : position = 8'd3;
        48'b00001??????????????????????????????????????????? : position = 8'd4;
        48'b000001?????????????????????????????????????????? : position = 8'd5;
        48'b0000001????????????????????????????????????????? : position = 8'd6;
        48'b00000001???????????????????????????????????????? : position = 8'd7;
        48'b000000001??????????????????????????????????????? : position = 8'd8;
        48'b0000000001?????????????????????????????????????? : position = 8'd9;
        48'b00000000001????????????????????????????????????? : position = 8'd10;
        48'b000000000001???????????????????????????????????? : position = 8'd11;
        48'b0000000000001??????????????????????????????????? : position = 8'd12;
        48'b00000000000001?????????????????????????????????? : position = 8'd13;
        48'b000000000000001????????????????????????????????? : position = 8'd14;
        48'b0000000000000001???????????????????????????????? : position = 8'd15;
        48'b00000000000000001??????????????????????????????? : position = 8'd16;
        48'b000000000000000001?????????????????????????????? : position = 8'd17;
        48'b0000000000000000001????????????????????????????? : position = 8'd18;
        48'b00000000000000000001???????????????????????????? : position = 8'd19;
        48'b000000000000000000001??????????????????????????? : position = 8'd20;
        48'b0000000000000000000001?????????????????????????? : position = 8'd21;
        48'b00000000000000000000001????????????????????????? : position = 8'd22;
        48'b000000000000000000000001???????????????????????? : position = 8'd23;
        default: position = 8'd24; // Assume denormalized
    endcase
end

//// Normalize Mantissa and Exponent
always @(*) begin
    if (exception) begin
        normalized_mantissa = 24'b0;
        normalized_exponent = 8'b0;
    end else begin
        shifted_mantissa = mantissa_div_result << position;  
        normalized_mantissa = shifted_mantissa[47:25];  // Take upper 23 bits
        normalized_exponent = adjusted_exponent - position;  
    end
end

assign pos = position;

// Calculate the output sign
always @(*) begin
    sign_out = sign_num1 ^ sign_num2;
end

// Combine the final result
always @(*) begin
    div_result = (exception) ? 32'b0 : {sign_out, normalized_exponent, normalized_mantissa};
end

endmodule
